module simplified_sha256 #(parameter integer NUM_OF_WORDS = 20)(
 input logic  clk, reset_n, start,
 input logic  [15:0] message_addr, output_addr,
 output logic done, mem_clk, mem_we,
 output logic [15:0] mem_addr,
 output logic [31:0] mem_write_data,
 input logic [31:0] mem_read_data);

// FSM state variables 
enum logic [2:0] {IDLE, READ, BLOCK, COMPUTE, WRITE} state;

// NOTE : Below mentioned frame work is for reference purpose.
// Local variables might not be complete and you might have to add more variables
// or modify these variables. Code below is more as a reference.

// Local variables
logic [31:0] w[16];
logic [31:0] message[20];
//logic [31:0] dpsram[0:16383];
//logic   [31:0] s1, s0;
logic [31:0] wt;
logic [31:0] h0, h1, h2, h3, h4, h5, h6, h7;
logic [31:0] a, b, c, d, e, f, g, h;
logic [ 7:0] i, j, n;
logic [15:0] offset; // in word address
logic [ 7:0] num_blocks;
logic        cur_we;			// write enabler 
logic [15:0] cur_addr;
logic [31:0] cur_write_data;
logic [512:0] memory_block;
//logic [ 7:0] tstep;

int t;

// SHA256 K constants
parameter int k[0:63] = '{
   32'h428a2f98,32'h71374491,32'hb5c0fbcf,32'he9b5dba5,32'h3956c25b,32'h59f111f1,32'h923f82a4,32'hab1c5ed5,
   32'hd807aa98,32'h12835b01,32'h243185be,32'h550c7dc3,32'h72be5d74,32'h80deb1fe,32'h9bdc06a7,32'hc19bf174,
   32'he49b69c1,32'hefbe4786,32'h0fc19dc6,32'h240ca1cc,32'h2de92c6f,32'h4a7484aa,32'h5cb0a9dc,32'h76f988da,
   32'h983e5152,32'ha831c66d,32'hb00327c8,32'hbf597fc7,32'hc6e00bf3,32'hd5a79147,32'h06ca6351,32'h14292967,
   32'h27b70a85,32'h2e1b2138,32'h4d2c6dfc,32'h53380d13,32'h650a7354,32'h766a0abb,32'h81c2c92e,32'h92722c85,
   32'ha2bfe8a1,32'ha81a664b,32'hc24b8b70,32'hc76c51a3,32'hd192e819,32'hd6990624,32'hf40e3585,32'h106aa070,
   32'h19a4c116,32'h1e376c08,32'h2748774c,32'h34b0bcb5,32'h391c0cb3,32'h4ed8aa4a,32'h5b9cca4f,32'h682e6ff3,
   32'h748f82ee,32'h78a5636f,32'h84c87814,32'h8cc70208,32'h90befffa,32'ha4506ceb,32'hbef9a3f7,32'hc67178f2
};


assign num_blocks = determine_num_blocks(NUM_OF_WORDS); 
//assign tstep = (i - 1);

// Note : Function defined are for reference purpose. Feel free to add more functions or modify below.
// Function to determine number of blocks in memory to fetch
function logic [15:0] determine_num_blocks(input logic [31:0] size);

  // Student to add function implementation
  determine_num_blocks = ((size * 32) / 512) + 1;
  

endfunction


// SHA256 hash round
function logic [255:0] sha256_op(input logic [31:0] a, b, c, d, e, f, g, h, w,
                                 input logic [7:0] t);
    logic [31:0] S1, S0, ch, maj, t1, t2; // internal signals
	 begin
		 S1 = rightrotate(e, 6) ^ rightrotate(e, 11) ^ rightrotate(e, 25);
		 // Student to add remaning code below
		 ch = (e & f) ^ ((~e) & g);
		 t1 = h + S1 + ch + k[t] + w;
		 S0 = rightrotate(a, 2) ^ rightrotate(a, 13) ^ rightrotate(a, 22);
		 maj = (a & b) ^ (a & c) ^ (b & c);
		 t2 = S0 + maj;
		 sha256_op = {t1 + t2, a, b, c, d + t1, e, f, g};
	 end
endfunction
// wtnew
function logic [31:0] wtnew; 
	logic [31:0] s1, s0;
	s0 = rightrotate(w[1], 7) ^ rightrotate(w[1], 18) ^ (w[1] >> 3);
   s1 = rightrotate(w[14], 17) ^ rightrotate(w[14], 19) ^ (w[14] >> 10);
   wtnew = w[0] + s0 + w[9] + s1;
endfunction
/*
function logic [31:0] wtnew(logic[7:0] t);
 logic [31:0] s1, s0;
 s0 = rightrotate(w[t-15], 7) ^ rightrotate(w[t-15], 18) ^ (w[t-15] >> 3);
 s1 = rightrotate(w[t-2], 17) ^ rightrotate(w[t-2], 19) ^ (w[t-2] >> 10);
 wtnew = w[t-16] + s0 + w[t-7] + s1;
endfunction
*/
// Generate request to memory
// for reading from memory to get original message
// for writing final computed has value
assign mem_clk = clk;
assign mem_addr = cur_addr + offset;
assign mem_we = cur_we;
assign mem_write_data = cur_write_data;


// Right Rotation Example : right rotate input x by r
// Lets say input x = 1111 ffff 2222 3333 4444 6666 7777 8888
// lets say r = 4
// x >> r  will result in : 0000 1111 ffff 2222 3333 4444 6666 7777 
// x << (32-r) will result in : 8888 0000 0000 0000 0000 0000 0000 0000
// final right rotate expression is = (x >> r) | (x << (32-r));
// (0000 1111 ffff 2222 3333 4444 6666 7777) | (8888 0000 0000 0000 0000 0000 0000 0000)
// final value after right rotate = 8888 1111 ffff 2222 3333 4444 6666 7777
// Right rotation function
function logic [31:0] rightrotate(input logic [31:0] x,
                                  input logic [ 7:0] r);
   // Student to add function implementation
	rightrotate = (x >> r) | (x << (32 - r));

endfunction


// SHA-256 FSM 
// Get a BLOCK from the memory, COMPUTE Hash output using SHA256 function
// and write back hash value back to memory
always_ff @(posedge clk, negedge reset_n)
begin
  if (!reset_n) begin
    cur_we <= 1'b0;
    state <= IDLE;
    offset <= 0;
  end 
 else case (state)
    IDLE: begin 
       if(start) begin
          //Initialize hash values:
          //(first 32 bits of the fractional parts of the square roots of the first 8 primes 2..19):
          h0 <= 32'h6a09e667;
          h1 <= 32'hbb67ae85;
          h2 <= 32'h3c6ef372;
          h3 <= 32'ha54ff53a;
          h4 <= 32'h510e527f;
          h5 <= 32'h9b05688c;
          h6 <= 32'h1f83d9ab;
          h7 <= 32'h5be0cd19;
	 
			 a <= 32'h0;
          b <= 32'h0;
          c <= 32'h0;
          d <= 32'h0;
          e <= 32'h0;
          f <= 32'h0;
          g <= 32'h0;
          h <= 32'h0;

          // Number of block iteration variable
          j <= 0;
     	    i <= 0;
			 
          // initialize pointer to access memory location
          offset <= 0;
	 
			 // by default set write enable to '0' (i.e. memory read mode)
          cur_we <= 1'b0;
			 
          // get starting address of message 
          cur_addr <= message_addr;
			 
			 // initialize write data to memory to '0'
          cur_write_data <= 32'h0;
			 
			 // proceed to message block fetch stage
			 state <= READ;
        end
    end
   
    // Read all input message words and store in vector array 'w'
    READ: begin
      if(offset<=20) begin
        if(offset != 0) begin
          message[offset-1] <= mem_read_data;
        end
      
       // Increment memory address to fetch next block 
       offset <= offset + 1;

       // stay in read memory state until all input message words are read
       state <= READ;
      end
      else begin
			offset <= 0;
         state <= BLOCK;
      end
    end	 

    // Create Both Blocks
    BLOCK: begin
		//i <= 0;
		if (j < num_blocks) begin
			if (j == 0) begin
				a <= h0;
				b <= h1;
				c <= h2;
				d <= h3;
				e <= h4;
				f <= h5;
				g <= h6;
				h <= h7;
				for (n = 0; n < 16; n++) w[n] <= message[n];
				
			end
			else begin
				a <= h0;
				b <= h1;
				c <= h2;
				d <= h3;
				e <= h4;
				f <= h5;
				g <= h6;
				h <= h7;
				
				for (n = 16; n < 20; n++) w[n-16] <= message[n];
				w[4] <= 32'h80000000;
				for (n = 21; n < 31; n++) w[n-16] <= 0;
				w[15] <= 32'd640;
			end
			state <= COMPUTE;
         i <= 0;
		end
		else begin
			i <= 0;
			state <= WRITE;
		end
   end

   // Perform word expansion and SHA256 operation
   COMPUTE: begin
       if (i <= 64) begin
          if(i<16) begin 
            {a,b,c,d,e,f,g,h} <= sha256_op(a, b, c, d, e, f, g, h, w[i], i);
          end
          else begin
				for (n = 0; n < 15; n++) w[n] <= w[n+1];
            w[15] <= wtnew(); // perform word expansion 
            // Since wtnew above mentioned line is non-blocking, the expanded w[16] to w[64] would take
            // 1 additional cycle to get its value available. Hence below mentioned guarded i!=16 in if block
            // where we do not do any SHA operation for 16th iteration as we are waiting for 1 cycle. From 17th iteration cycle
            // we perform SHA operation. Also note that due to this 1 dummy cycle of not doing anything when 
            // i moves to 17, then w[i-1] and i-1 are used in sha256_op below to compute SHA operation for w[16] word
            // And hence i<=64 used in above mentioned if(i<=64) line insted of if(i<64)
            if(i != 16) {a,b,c,d,e,f,g,h} <= sha256_op(a, b, c, d, e, f, g, h, w[15], i-1);
          end
          i <= i + 1;
			 state <= COMPUTE;
       end
       else begin
			 h0 <= h0 + a;
			 h1 <= h1 + b;
			 h2 <= h2 + c;
			 h3 <= h3 + d;
			 h4 <= h4 + e;
			 h5 <= h5 + f;
			 h6 <= h6 + g;
			 h7 <= h7 + h;
			 state <= BLOCK;
			 j <= j + 1;
		 end
    end

    // Write output hash value back to the memory
    WRITE: begin
		if (i <= 7) begin 
			state <= WRITE;
			i <= i + 1;
			offset <= i;
			cur_we <= 1'b1;
         cur_addr <= output_addr;
			if (i == 0)
				cur_write_data <= h0;
			else if (i == 1)
				cur_write_data <= h1;
			else if (i == 2) 
				cur_write_data <= h2;
			else if (i == 3) 
				cur_write_data <= h3;
			else if (i == 4) 
				cur_write_data <= h4;
			else if (i == 5)
				cur_write_data <= h5;
			else if (i == 6)
				cur_write_data <= h6;
			else if (i == 7)
				cur_write_data <= h7;
		end
		else begin
			cur_we <= 1'b0;
			offset <= 0;
			state <= IDLE;
			i <= 0;
		end	
    end
   endcase
end


// Generate done when SHA256 hash computation has finished and moved to IDLE state
assign done = (state == IDLE);

endmodule




